

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_top is

end tb_top;

architecture testbench of tb_top is
    component top
        Port ( 
            clk: in std_logic;
            reset: in std_logic;
            speed: in std_logic;
            mode: in std_logic_vector (1 downto 0);
            B4: in std_logic;
            B3: in std_logic;
            B2: in std_logic;
            B1: in std_logic;
            selector: out std_logic_vector (3 downto 0);
            segmentos: out std_logic_vector (7 downto 0);
            leds: out std_logic_vector (7 downto 0)
            );
    end component;
    
    signal clk: std_logic;
    signal reset: std_logic;
    signal speed: std_logic;
    signal mode: std_logic_vector (1 downto 0);
    signal B4: std_logic;
    signal B3: std_logic;
    signal B2: std_logic;
    signal B1: std_logic;
    signal selector: std_logic_vector (3 downto 0);
    signal segmentos: std_logic_vector (7 downto 0);
    signal leds: std_logic_vector (7 downto 0);
    
    
    --declaracion tiempo
    constant clk_period_real : time := 8 ns;
    constant clk_period : time := 800ns;

    begin
    
    --instanciacion componente
    uut: top
    port map (
        clk => clk,
        reset => reset,
        speed => speed,
        mode => mode,
        B4 => B4,
        B3 => B3,
        B2 => B2,
        B1 => B1,
        selector => selector,
        segmentos => segmentos,
        leds => leds
    );
    
     --generacion de reloj
     process
     begin
         clk <= '1';
         wait for clk_period_real/2;
         clk <= '0';
         wait for clk_period_real/2;        
     end process;
     
     --generacion resto de entradas
     process
     begin
         reset <= '1';
         speed <= '1';
         mode <= "00";
         B4 <= '0';
         B3 <= '0';
         B2 <= '0';
         B1 <= '0';
        
         wait for clk_period*200;
         reset <= '0';
         wait for clk_period*100;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0';
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0'; 
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*2000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';   
         wait for clk_period*100;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         
                  
         
         wait for clk_period*10000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*2000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';   
         
         
         wait for clk_period*20000;
         reset <= '0';
         wait for clk_period*100;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0';
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0'; 
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B2 <= '1';
         wait for clk_period*2000;
         B2 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*2000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';   
         wait for clk_period*100;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         
                  
         
         wait for clk_period*10000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*2000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         
                  wait for clk_period*20000;
         reset <= '0';
         wait for clk_period*100;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0';
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0'; 
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B2 <= '1';
         wait for clk_period*2000;
         B2 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*2000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';   
         wait for clk_period*100;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         
                  
         
         wait for clk_period*10000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*2000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         
                  wait for clk_period*20000;
         reset <= '0';
         wait for clk_period*100;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0';
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0'; 
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B2 <= '1';
         wait for clk_period*2000;
         B2 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*2000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';   
         wait for clk_period*100;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         
                  
         
         wait for clk_period*10000;
         B2 <= '1';
         wait for clk_period*500;
         B2 <= '0';
         wait for clk_period*100;
         B1 <= '1';
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B3 <= '1';
         wait for clk_period*500;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B4 <= '1';
         wait for clk_period*500;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*1000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*1000;
         B4 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait for clk_period*1000;
         B3 <= '1';
         wait for clk_period*1000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';  
         wait for clk_period*500;
         B2 <= '1';
         wait for clk_period*2000;
         B2 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';                             
         wait for clk_period*1000;
         B4 <= '1';
         wait for clk_period*2000;
         B4 <= '0'; 
         wait for clk_period*500;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';    
         wait for clk_period*2000;
         B3 <= '1';
         wait for clk_period*2000;
         B3 <= '0'; 
         wait for clk_period*1000;
         B1 <= '1';  
         wait for clk_period*1000;
         B1 <= '0';
         wait;
    end process;
       
end testbench;
